*Ejemplo de plataforma de entrada de SPICE para un 
*circuito simple divisor de tensión.

R1 1 2 1k
R2 2 0 1k
V1 1 0 5
*Solicita el punto de operación de DC
.op
.end